
module MyAnd (
 input a,
 input b,
 output c
);
 
 // Puerta and
 
 assign 
 c=a&b;
 
endmodule
