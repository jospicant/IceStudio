
module triestadop(inout pin,input in,input eo);

bufif1 myBufferP(pin,in,eo);

endmodule
