
module MyAnd (
 input a,
 input b,
 output o
);
 
 //AND
 
 assign o=a&b;
endmodule
