
module triestadon(inout pin,input in,input eo);

bufif0 myBufferN(pin,in,eo);

endmodule
