
//En función de si comento o no EleccionA tendré un resultado u otro 

`define EleccionA

`define A 4'b0101
`define B 4'b1010
